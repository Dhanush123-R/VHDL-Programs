LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FULLSUB IS
PORT(
A,BIN,C : IN STD_LOGIC;
D,BOUT : OUT STD_LOGIC
);
END FULLSUB;

ARCHITECTURE DATAFLOW OF FULLSUB IS
BEGIN
D <= A XOR BIN XOR C;
BOUT <= ((BIN XOR C) AND (NOT A)) OR (BIN AND C);
END DATAFLOW;
